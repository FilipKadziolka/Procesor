//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "procesor.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
wire w6;    //: /sn:0 {0}(735,222)(735,237){1}
wire w32;    //: /sn:0 {0}(708,408)(708,423){1}
wire w7;    //: /sn:0 {0}(700,222)(700,237){1}
wire w45;    //: /sn:0 {0}(339,408)(339,423){1}
wire w46;    //: /sn:0 {0}(321,408)(321,423){1}
wire w14;    //: /sn:0 {0}(539,211)(539,226){1}
wire w16;    //: /sn:0 {0}(435,124)(435,109){1}
wire w56;    //: /sn:0 {0}(306,481)(306,466){1}
wire w4;    //: /sn:0 {0}(731,129)(731,114){1}
wire w15;    //: /sn:0 {0}(504,211)(504,226){1}
wire w19;    //: /sn:0 {0}(404,217)(404,232){1}
wire w38;    //: /sn:0 {0}(594,408)(594,423){1}
wire w51;    //: /sn:0 {0}(510,481)(510,466){1}
wire w3;    //: /sn:0 {0}(827,224)(827,209){1}
wire w0;    //: /sn:0 {0}(787,101)(787,116){1}
wire w37;    //: /sn:0 {0}(612,408)(612,423){1}
wire w34;    //: /sn:0 {0}(667,408)(667,423){1}
wire w21;    //: /sn:0 {0}(314,128)(314,113){1}
wire w43;    //: /sn:0 {0}(375,408)(375,423){1}
wire w54;    //: /sn:0 {0}(448,481)(448,466){1}
wire w31;    //: /sn:0 {0}(120,230)(120,245){1}
wire w28;    //: /sn:0 {0}(151,137)(151,122){1}
wire w20;    //: /sn:0 {0}(350,128)(350,113){1}
wire w23;    //: /sn:0 {0}(319,221)(319,236){1}
wire w24;    //: /sn:0 {0}(245,127)(245,112){1}
wire w36;    //: /sn:0 {0}(629,408)(629,423){1}
wire w41;    //: /sn:0 {0}(410,408)(410,423){1}
wire w1;    //: /sn:0 {0}(823,101)(823,116){1}
wire w25;    //: /sn:0 {0}(209,127)(209,112){1}
wire w8;    //: /sn:0 {0}(618,118)(618,103){1}
wire w18;    //: /sn:0 {0}(439,217)(439,232){1}
wire w35;    //: /sn:0 {0}(650,408)(650,423){1}
wire w40;    //: /sn:0 {0}(424,408)(424,423){1}
wire w30;    //: /sn:0 {0}(155,230)(155,245){1}
wire w17;    //: /sn:0 {0}(399,124)(399,109){1}
wire w22;    //: /sn:0 {0}(354,221)(354,236){1}
wire w53;    //: /sn:0 {0}(467,481)(467,466){1}
wire w2;    //: /sn:0 {0}(792,224)(792,209){1}
wire w11;    //: /sn:0 {0}(587,211)(587,226){1}
wire w12;    //: /sn:0 {0}(535,118)(535,103){1}
wire w44;    //: /sn:0 {0}(359,408)(359,423){1}
wire w49;    //: /sn:0 {0}(559,481)(559,466){1}
wire w10;    //: /sn:0 {0}(622,211)(622,226){1}
wire w13;    //: /sn:0 {0}(499,118)(499,103){1}
wire w27;    //: /sn:0 {0}(214,220)(214,235){1}
wire w5;    //: /sn:0 {0}(695,129)(695,114){1}
wire w33;    //: /sn:0 {0}(688,408)(688,423){1}
wire w48;    //: /sn:0 {0}(585,481)(585,466){1}
wire w52;    //: /sn:0 {0}(485,481)(485,466){1}
wire w29;    //: /sn:0 {0}(115,137)(115,122){1}
wire w47;    //: /sn:0 {0}(296,408)(296,423){1}
wire w9;    //: /sn:0 {0}(582,118)(582,103){1}
wire w42;    //: /sn:0 {0}(394,408)(394,423){1}
wire w50;    //: /sn:0 {0}(535,481)(535,466){1}
wire w26;    //: /sn:0 {0}(249,220)(249,235){1}
wire w39;    //: /sn:0 {0}(574,408)(574,423){1}
wire w55;    //: /sn:0 {0}(426,481)(426,466){1}
//: enddecls

  generacja g4 (.x(w17), .y(w16), .g(w19), .h(w18));   //: @(380, 125) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  sumator g8 (.y7(w47), .y6(w46), .y5(w45), .y4(w44), .y3(w43), .y2(w42), .y1(w41), .y0(w40), .x7(w39), .x6(w38), .x5(w37), .x4(w36), .x3(w35), .x2(w34), .x1(w33), .x0(w32), .c8(w56), .s7(w55), .s6(w54), .s5(w53), .s4(w52), .s3(w51), .s2(w50), .s1(w49), .s0(w48));   //: @(237, 424) /sz:(500, 41) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ti8>1 Ti9>1 Ti10>1 Ti11>1 Ti12>1 Ti13>1 Ti14>1 Ti15>1 Bo0<1 Bo1<1 Bo2<1 Bo3<1 Bo4<1 Bo5<1 Bo6<1 Bo7<1 Bo8<1 ]
  generacja g3 (.x(w13), .y(w12), .g(w15), .h(w14));   //: @(480, 119) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g2 (.x(w9), .y(w8), .g(w11), .h(w10));   //: @(563, 119) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g1 (.x(w5), .y(w4), .g(w7), .h(w6));   //: @(676, 130) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g6 (.x(w25), .y(w24), .g(w27), .h(w26));   //: @(190, 128) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g7 (.x(w29), .y(w28), .g(w31), .h(w30));   //: @(96, 138) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g5 (.x(w21), .y(w20), .g(w23), .h(w22));   //: @(295, 129) /sz:(82, 91) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Bo1<0 ]
  generacja g0 (.y(w1), .x(w0), .h(w3), .g(w2));   //: @(768, 117) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin generacja
module generacja(y, h, g, x);
//: interface  /sz:(82, 91) /bd:[ Ti0>x(19/82) Ti1>y(55/82) Bo0<g(24/82) Bo1<h(59/82) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output h;    //: /sn:0 {0}(401,296)(401,259){1}
input y;    //: /sn:0 {0}(405,156)(405,191)(405,191)(405,194){1}
//: {2}(403,196)(346,196)(346,235){3}
//: {4}(405,198)(405,225)(404,225)(404,238){5}
input x;    //: /sn:0 {0}(333,152)(333,178){1}
//: {2}(335,180)(399,180)(399,238){3}
//: {4}(333,182)(333,222)(341,222)(341,235){5}
output g;    //: /sn:0 {0}(343,256)(343,310){1}
//: enddecls

  //: joint g4 (y) @(405, 196) /w:[ -1 1 2 4 ]
  _GGXOR2 #(8) g3 (.I0(y), .I1(x), .Z(h));   //: @(401,249) /sn:0 /R:3 /w:[ 5 3 1 ]
  _GGAND2 #(6) g2 (.I0(y), .I1(x), .Z(g));   //: @(343,246) /sn:0 /R:3 /w:[ 3 5 0 ]
  //: IN g1 (y) @(405,154) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g6 (h) @(401,293) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g7 (g) @(343,307) /sn:0 /R:3 /w:[ 1 ]
  //: joint g5 (x) @(333, 180) /w:[ 2 1 -1 4 ]
  //: IN g0 (x) @(333,150) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin sumator
module sumator();
//: interface  /sz:(500, 41) /bd:[ Ti0>y7(59/500) Ti1>y6(84/500) Ti2>y5(102/500) Ti3>y4(122/500) Ti4>y3(138/500) Ti5>y2(157/500) Ti6>y1(173/500) Ti7>y0(187/500) Ti8>x7(337/500) Ti9>x6(357/500) Ti10>x5(375/500) Ti11>x4(392/500) Ti12>x3(413/500) Ti13>x2(430/500) Ti14>x1(451/500) Ti15>x0(471/500) Bo0<c8(69/500) Bo1<s7(189/500) Bo2<s6(211/500) Bo3<s5(230/500) Bo4<s4(248/500) Bo5<s3(273/500) Bo6<s2(298/500) Bo7<s1(322/500) Bo8<s0(348/500) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
//: enddecls


endmodule
//: /netlistEnd

