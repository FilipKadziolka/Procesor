//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "procesor.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w6;    //: /sn:0 {0}(594,423)(594,396)(565,396)(565,324){1}
reg w7;    //: /sn:0 {0}(536,287)(536,408)(574,408)(574,423){1}
reg w14;    //: /sn:0 {0}(321,423)(321,394)(296,394)(296,318){1}
reg w15;    //: /sn:0 {0}(265,284)(265,403)(296,403)(296,423){1}
reg w4;    //: /sn:0 {0}(623,324)(623,408)(0:629,408)(629,423){1}
reg w0;    //: /sn:0 {0}(708,423)(708,408)(738,408)(738,325){1}
reg w3;    //: /sn:0 {0}(648,290)(648,408)(650,408)(650,423){1}
reg w1;    //: /sn:0 {0}(688,423)(688,399)(707,399)(707,290){1}
reg w8;    //: /sn:0 {0}(443,316)(443,408)(424,408)(424,423){1}
reg w12;    //: /sn:0 {0}(359,423)(359,393)(343,393)(343,320){1}
reg w11;    //: /sn:0 {0}(375,423)(375,394)(369,394)(369,286){1}
reg w2;    //: /sn:0 {0}(677,324)(677,408)(667,408)(667,423){1}
reg w10;    //: /sn:0 {0}(393,321)(393,408)(394,408)(394,423){1}
reg w13;    //: /sn:0 {0}(339,423)(339,387)(322,387)(322,279){1}
reg w5;    //: /sn:0 {0}(612,423)(612,390)(591,390)(591,284){1}
reg w9;    //: /sn:0 {0}(410,423)(410,390)(421,390)(421,285){1}
wire w56;    //: /sn:0 {0}(306,466)(306,499)(307,499)(307,514){1}
wire w51;    //: /sn:0 {0}(510,466)(510,497)(511,497)(511,512){1}
wire w54;    //: /sn:0 {0}(448,466)(448,488)(451,488)(451,510){1}
wire w53;    //: /sn:0 {0}(467,466)(467,506){1}
wire w49;    //: /sn:0 {0}(559,466)(559,517){1}
wire w48;    //: /sn:0 {0}(585,466)(585,508)(587,508)(587,523){1}
wire w52;    //: /sn:0 {0}(485,466)(485,499)(488,499)(488,514){1}
wire w50;    //: /sn:0 {0}(535,466)(535,516){1}
wire w55;    //: /sn:0 {0}(427,504)(427,481)(426,481)(426,466){1}
//: enddecls

  sumator g8 (.y7(w15), .y6(w14), .y5(w13), .y4(w12), .y3(w11), .y2(w10), .y1(w9), .y0(w8), .x7(w7), .x6(w6), .x5(w5), .x4(w4), .x3(w3), .x2(w2), .x1(w1), .x0(w0), .c8(w56), .s7(w55), .s6(w54), .s5(w53), .s4(w52), .s3(w51), .s2(w50), .s1(w49), .s0(w48));   //: @(237, 424) /sz:(500, 41) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>1 Ti6>0 Ti7>1 Ti8>1 Ti9>0 Ti10>0 Ti11>1 Ti12>1 Ti13>1 Ti14>0 Ti15>0 Bo0<0 Bo1<1 Bo2<0 Bo3<0 Bo4<0 Bo5<0 Bo6<0 Bo7<0 Bo8<0 ]
  //: SWITCH g4 (w4) @(623,311) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g13 (w12) @(343,307) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g3 (w3) @(648,277) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g2 (w2) @(677,311) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g1 (w1) @(707,277) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g16 (w15) @(265,271) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g11 (w10) @(393,308) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g10 (w9) @(421,272) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: LED g19 (w50) @(535,523) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g6 (w6) @(565,311) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g7 (w7) @(536,274) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g9 (w8) @(443,303) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: LED g20 (w51) @(511,519) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g15 (w14) @(296,305) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: LED g25 (w56) @(307,521) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: LED g17 (w48) @(587,530) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g14 (w13) @(322,266) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g5 (w5) @(591,271) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: LED g24 (w55) @(427,511) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: LED g21 (w52) @(488,521) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: LED g23 (w54) @(451,517) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: LED g22 (w53) @(467,513) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g0 (w0) @(738,312) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1
  //: LED g18 (w49) @(559,524) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g12 (w11) @(369,273) /sn:0 /R:3 /w:[ 1 ] /st:0 /dn:1

endmodule
//: /netlistEnd

//: /netlistBegin generacja
module generacja(y, h, g, x);
//: interface  /sz:(82, 91) /bd:[ Ti0>x(19/82) Ti1>y(55/82) Bo0<g(24/82) Bo1<h(59/82) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output h;    //: /sn:0 {0}(401,296)(401,259){1}
input y;    //: /sn:0 {0}(405,156)(405,191)(405,191)(405,194){1}
//: {2}(403,196)(346,196)(346,235){3}
//: {4}(405,198)(405,225)(404,225)(404,238){5}
input x;    //: /sn:0 {0}(333,152)(333,178){1}
//: {2}(335,180)(399,180)(399,238){3}
//: {4}(333,182)(333,222)(341,222)(341,235){5}
output g;    //: /sn:0 {0}(343,256)(343,310){1}
//: enddecls

  //: joint g4 (y) @(405, 196) /w:[ -1 1 2 4 ]
  _GGXOR2 #(8) g3 (.I0(y), .I1(x), .Z(h));   //: @(401,249) /sn:0 /R:3 /w:[ 5 3 1 ]
  _GGAND2 #(6) g2 (.I0(y), .I1(x), .Z(g));   //: @(343,246) /sn:0 /R:3 /w:[ 3 5 0 ]
  //: IN g1 (y) @(405,154) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g6 (h) @(401,293) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g7 (g) @(343,307) /sn:0 /R:3 /w:[ 1 ]
  //: joint g5 (x) @(333, 180) /w:[ 2 1 -1 4 ]
  //: IN g0 (x) @(333,150) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin sumator
module sumator(y0, s3, y5, c8, s4, x0, y3, s6, y2, x3, s1, y1, x4, y7, s5, x1, y6, x5, s7, s2, x7, x6, x2, y4, s0);
//: interface  /sz:(500, 41) /bd:[ Ti0>y7(59/500) Ti1>y6(84/500) Ti2>y5(102/500) Ti3>y4(122/500) Ti4>y3(138/500) Ti5>y2(157/500) Ti6>y1(173/500) Ti7>y0(187/500) Ti8>x7(337/500) Ti9>x6(357/500) Ti10>x5(375/500) Ti11>x4(392/500) Ti12>x3(413/500) Ti13>x2(430/500) Ti14>x1(451/500) Ti15>x0(471/500) Bo0<c8(69/500) Bo1<s7(189/500) Bo2<s6(211/500) Bo3<s5(230/500) Bo4<s4(248/500) Bo5<s3(273/500) Bo6<s2(298/500) Bo7<s1(322/500) Bo8<s0(348/500) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output s2;    //: /sn:0 {0}(656,696)(656,644)(650,644)(650,629){1}
input x1;    //: /sn:0 {0}(663,32)(663,47)(669,47)(669,77){1}
output s0;    //: /sn:0 {0}(799,170)(799,289){1}
//: {2}(801,291)(809,291)(809,623){3}
//: {4}(797,291)(722,291)(722,306){5}
input y4;    //: /sn:0 {0}(412,30)(412,50)(413,50)(413,77){1}
output s6;    //: /sn:0 {0}(248,750)(248,810){1}
input x0;    //: /sn:0 {0}(755,32)(755,50)(759,50)(759,77){1}
output c8;    //: /sn:0 {0}(7,757)(7,794)(6,794)(6,809){1}
input y0;    //: /sn:0 {0}(799,32)(799,59)(795,59)(795,77){1}
input x7;    //: /sn:0 {0}(102,29)(102,55)(100,55)(100,77){1}
output s3;    //: /sn:0 {0}(591,521)(591,615)(594,615)(594,675){1}
output s1;    //: /sn:0 {0}(762,613)(762,651)(763,651)(763,666){1}
input x4;    //: /sn:0 {0}(372,32)(372,63)(377,63)(377,77){1}
output s4;    //: /sn:0 {0}(457,714)(457,759)(462,759)(462,763){1}
input y1;    //: /sn:0 {0}(703,32)(703,54)(705,54)(705,77){1}
input y2;    //: /sn:0 {0}(610,32)(610,35)(609,35)(609,43){1}
//: {2}(611,45)(617,45){3}
//: {4}(609,47)(609,77){5}
input x6;    //: /sn:0 {0}(203,33)(203,55)(201,55)(201,77){1}
output s5;    //: /sn:0 {0}(377,736)(377,782)(382,782)(382,792){1}
input x3;    //: /sn:0 {0}(462,32)(462,66)(468,66)(468,77){1}
input y3;    //: /sn:0 {0}(504,63)(504,66){1}
//: {2}(502,68)(492,68)(492,51)(506,51)(506,34){3}
//: {4}(504,70)(504,77){5}
input x5;    //: /sn:0 {0}(294,31)(294,49)(288,49){1}
//: {2}(286,47)(286,42){3}
//: {4}(286,51)(286,53)(290,53)(290,77){5}
output s7;    //: /sn:0 {0}(156,744)(156,801)(160,801)(160,808){1}
input y5;    //: /sn:0 {0}(325,31)(325,66)(326,66)(326,77){1}
input y7;    //: /sn:0 {0}(136,30)(136,77){1}
input x2;    //: /sn:0 {0}(564,32)(564,49)(573,49)(573,77){1}
input y6;    //: /sn:0 {0}(235,31)(235,61)(237,61)(237,77){1}
wire w32;    //: /sn:0 {0}(-7,692)(-7,592)(26,592)(26,541){1}
wire w6;    //: /sn:0 {0}(674,170)(674,226)(654,226)(654,253)(655,253)(655,263){1}
//: {2}(653,265)(647,265){3}
//: {4}(655,267)(655,277)(646,277)(646,306){5}
wire w7;    //: /sn:0 {0}(709,170)(709,248){1}
//: {2}(711,250)(760,250)(760,592){3}
//: {4}(707,250)(681,250)(681,264)(678,264){5}
//: {6}(674,264)(668,264){7}
//: {8}(676,266)(676,276)(663,276)(663,306){9}
wire w16;    //: /sn:0 {0}(71,476)(71,461)(50,461)(50,449)(155,449){1}
//: {2}(159,449)(248,449){3}
//: {4}(252,449)(267,449)(267,370){5}
//: {6}(250,451)(250,474)(244,474)(244,498){7}
//: {8}(157,451)(157,472)(155,472)(155,482){9}
wire w14;    //: /sn:0 {0}(450,295)(450,259)(473,259)(473,170){1}
wire w4;    //: /sn:0 {0}(124,305)(124,285)(239,285){1}
//: {2}(241,283)(241,170){3}
//: {4}(241,287)(241,295)(231,295)(231,391)(239,391)(239,471){5}
//: {6}(237,473)(221,473)(221,497){7}
//: {8}(239,475)(239,498){9}
wire w19;    //: /sn:0 {0}(417,170)(417,289){1}
//: {2}(415,291)(329,291)(329,305){3}
//: {4}(417,293)(417,599)(455,599)(455,663){5}
//: {6}(453,665)(400,665)(400,688){7}
//: {8}(455,667)(455,693){9}
wire w15;    //: /sn:0 {0}(508,170)(508,246){1}
//: {2}(510,248)(565,248)(565,350){3}
//: {4}(508,250)(508,271)(467,271)(467,295){5}
wire w38;    //: /sn:0 {0}(104,452)(104,458){1}
//: {2}(106,460)(176,460){3}
//: {4}(180,460)(211,460){5}
//: {6}(215,460)(270,460){7}
//: {8}(274,460)(296,460)(296,370){9}
//: {10}(272,462)(272,472)(271,472)(271,702){11}
//: {12}(213,462)(213,472)(216,472)(216,497){13}
//: {14}(178,462)(178,472)(175,472)(175,482){15}
//: {16}(104,462)(104,470)(88,470)(88,476){17}
wire w3;    //: /sn:0 {0}(567,371)(567,458)(575,458)(575,473){1}
wire w21;    //: /sn:0 {0}(660,371)(660,405){1}
//: {2}(658,407)(614,407){3}
//: {4}(610,407)(596,407){5}
//: {6}(592,407)(511,407)(511,521){7}
//: {8}(594,409)(594,473){9}
//: {10}(612,409)(612,419)(614,419)(614,473){11}
//: {12}(660,409)(660,595)(653,595)(653,608){13}
wire w31;    //: /sn:0 {0}(140,170)(140,238){1}
//: {2}(142,240)(159,240)(159,334){3}
//: {4}(140,242)(140,245)(65,245)(65,305){5}
wire w28;    //: /sn:0 {0}(36,757)(36,772){1}
wire w36;    //: /sn:0 {0}(136,482)(136,435)(161,435)(161,355){1}
wire w24;    //: /sn:0 {0}(537,444)(550,444){1}
//: {2}(554,444)(689,444)(689,371){3}
//: {4}(552,442)(552,440)(545,440)(545,446)(528,446)(528,521){5}
wire w20;    //: /sn:0 {0}(469,521)(469,488)(493,488)(493,360){1}
wire w23;    //: /sn:0 {0}(270,305)(270,275)(330,275)(330,262){1}
//: {2}(332,260)(367,260)(367,342){3}
//: {4}(330,258)(330,170){5}
wire w25;    //: /sn:0 {0}(69,692)(69,659)(92,659)(92,649){1}
//: {2}(94,647)(458,647){3}
//: {4}(462,647)(495,647)(495,586){5}
//: {6}(460,649)(460,693){7}
//: {8}(90,647)(84,647){9}
wire w35;    //: /sn:0 {0}(218,518)(218,681)(179,681)(179,696){1}
wire w8;    //: /sn:0 {0}(33,425)(39,425){1}
//: {2}(43,425)(62,425)(62,370){3}
//: {4}(41,423)(41,420)(12,420)(12,476){5}
wire w18;    //: /sn:0 {0}(382,170)(382,283)(373,283){1}
//: {2}(369,283)(312,283)(312,305){3}
//: {4}(371,285)(371,295)(372,295)(372,342){5}
wire w30;    //: /sn:0 {0}(105,170)(105,239)(48,239)(48,305){1}
wire w22;    //: /sn:0 {0}(295,170)(295,265)(253,265)(253,305){1}
wire w12;    //: /sn:0 {0}(52,692)(52,638)(63,638)(63,628){1}
//: {2}(65,626)(159,626){3}
//: {4}(163,626)(247,626){5}
//: {6}(251,626)(376,626){7}
//: {8}(380,626)(466,626)(466,586){9}
//: {10}(378,628)(378,640)(380,640)(380,688){11}
//: {12}(249,628)(249,638)(251,638)(251,702){13}
//: {14}(161,628)(161,638)(159,638)(159,696){15}
//: {16}(61,626)(52,626){17}
wire w11;    //: /sn:0 {0}(613,170)(613,278){1}
//: {2}(611,280)(526,280)(526,295){3}
//: {4}(613,282)(613,378)(648,378)(648,608){5}
wire w2;    //: /sn:0 {0}(705,306)(705,274)(762,274){1}
//: {2}(764,272)(764,170){3}
//: {4}(764,276)(764,472)(765,472)(765,592){5}
wire w10;    //: /sn:0 {0}(578,170)(578,266)(573,266){1}
//: {2}(569,266)(516,266)(516,272)(509,272)(509,295){3}
//: {4}(571,268)(571,278)(570,278)(570,350){5}
wire w27;    //: /sn:0 {0}(241,519)(241,687)(232,687)(232,702){1}
wire w13;    //: /sn:0 {0}(464,360)(464,481)(452,481)(452,521){1}
wire w33;    //: /sn:0 {0}(10,692)(10,621)(22,621)(22,611){1}
//: {2}(24,609)(55,609)(55,541){3}
//: {4}(20,609)(14,609){5}
wire w29;    //: /sn:0 {0}(369,363)(369,673)(361,673)(361,688){1}
wire w9;    //: /sn:0 {0}(91,370)(91,440)(29,440)(29,476){1}
wire w39;    //: /sn:0 {0}(140,696)(140,550)(152,550)(152,530){1}
wire w26;    //: /sn:0 {0}(107,305)(107,268)(163,268){1}
//: {2}(167,268)(206,268)(206,170){3}
//: {4}(165,270)(165,274)(164,274)(164,334){5}
//: enddecls

  _GGXOR2 #(8) g61 (.I0(w25), .I1(w19), .Z(s4));   //: @(457,704) /sn:0 /R:3 /w:[ 7 9 0 ]
  //: IN g8 (y0) @(799,30) /sn:0 /R:3 /w:[ 0 ]
  generacja g4 (.y(y4), .x(x4), .h(w19), .g(w18));   //: @(358, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  modul1 g58 (.Pi(w38), .Gi(w16), .Pk(w9), .Gk(w8), .Pki(w33), .Gki(w32));   //: @(-4, 477) /sz:(107, 63) /sn:0 /p:[ Ti0>17 Ti1>0 Ti2>1 Ti3>5 Bo0<3 Bo1<1 ]
  //: joint g55 (w18) @(371, 283) /w:[ 1 -1 2 4 ]
  //: OUT g51 (s3) @(594,672) /sn:0 /R:3 /w:[ 1 ]
  //: joint g37 (w7) @(709, 250) /w:[ 2 1 4 -1 ]
  //: joint g34 (s0) @(799, 291) /w:[ 2 1 4 -1 ]
  //: IN g13 (y5) @(325,29) /sn:0 /R:3 /w:[ 0 ]
  generacja g3 (.y(y3), .x(x3), .h(w15), .g(w14));   //: @(449, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>5 Ti1>1 Bo0<0 Bo1<1 ]
  //: joint g86 (w12) @(63, 626) /w:[ 2 -1 16 1 ]
  //: OUT g89 (c8) @(6,806) /sn:0 /R:3 /w:[ 1 ]
  //: joint g77 (w12) @(249, 626) /w:[ 6 -1 5 12 ]
  //: joint g76 (w38) @(272, 460) /w:[ 8 -1 7 10 ]
  modul2 g65 (.H(w19), .G(w12), .S(w29), .Sk(s5));   //: @(349, 689) /sz:(60, 46) /sn:0 /p:[ Ti0>7 Ti1>11 Ti2>1 Bo0<0 ]
  generacja g2 (.y(y2), .x(x2), .h(w11), .g(w10));   //: @(554, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>5 Ti1>1 Bo0<0 Bo1<0 ]
  //: joint g59 (w8) @(41, 425) /w:[ 2 4 1 -1 ]
  //: joint g72 (w4) @(241, 285) /w:[ -1 2 1 4 ]
  generacja g1 (.y(y1), .x(x1), .h(w7), .g(w6));   //: @(650, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  //: OUT g64 (s4) @(462,760) /sn:0 /R:3 /w:[ 1 ]
  //: IN g16 (x0) @(755,30) /sn:0 /R:3 /w:[ 0 ]
  //: IN g11 (y3) @(506,32) /sn:0 /R:3 /w:[ 3 ]
  //: OUT g78 (s6) @(248,807) /sn:0 /R:3 /w:[ 1 ]
  //: joint g50 (w21) @(612, 407) /w:[ 3 -1 4 10 ]
  modul1 g28 (.Pi(w19), .Gi(w18), .Pk(w23), .Gk(w22), .Pki(w38), .Gki(w16));   //: @(237, 306) /sz:(107, 63) /sn:0 /p:[ Ti0>3 Ti1>3 Ti2>0 Ti3>1 Bo0<9 Bo1<5 ]
  //: IN g10 (y2) @(610,30) /sn:0 /R:3 /w:[ 0 ]
  //: joint g87 (w25) @(92, 647) /w:[ 2 -1 8 1 ]
  //: joint g32 (w7) @(676, 264) /w:[ 5 -1 6 8 ]
  modul1 g27 (.Pi(w4), .Gi(w26), .Pk(w31), .Gk(w30), .Pki(w9), .Gki(w8));   //: @(32, 306) /sz:(107, 63) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>5 Ti3>1 Bo0<0 Bo1<3 ]
  //: IN g19 (x3) @(462,30) /sn:0 /R:3 /w:[ 0 ]
  _GGXOR2 #(8) g69 (.I0(w16), .I1(w4), .Z(w27));   //: @(241,509) /sn:0 /R:3 /w:[ 7 9 0 ]
  //: OUT g38 (s1) @(763,663) /sn:0 /R:3 /w:[ 1 ]
  generacja g6 (.y(y6), .x(x6), .h(w4), .g(w26));   //: @(182, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<3 Bo1<3 ]
  modul2 g75 (.H(w38), .G(w12), .S(w27), .Sk(s6));   //: @(220, 703) /sz:(60, 46) /sn:0 /p:[ Ti0>11 Ti1>13 Ti2>1 Bo0<0 ]
  //: joint g57 (w26) @(165, 268) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g53 (.I0(w18), .I1(w23), .Z(w29));   //: @(369,353) /sn:0 /R:3 /w:[ 5 3 0 ]
  //: IN g9 (y1) @(703,30) /sn:0 /R:3 /w:[ 0 ]
  generacja g7 (.y(y7), .x(x7), .h(w31), .g(w30));   //: @(81, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  modul2 g71 (.H(w38), .G(w16), .S(w36), .Sk(w39));   //: @(124, 483) /sz:(60, 46) /sn:0 /p:[ Ti0>15 Ti1>9 Ti2>0 Bo0<1 ]
  //: joint g31 (w6) @(655, 265) /w:[ -1 1 2 4 ]
  //: IN g20 (x4) @(372,30) /sn:0 /R:3 /w:[ 0 ]
  //: IN g15 (y7) @(136,28) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g68 (s5) @(382,789) /sn:0 /R:3 /w:[ 1 ]
  //: joint g67 (w12) @(378, 626) /w:[ 8 -1 7 10 ]
  _GGXOR2 #(8) g39 (.I0(w21), .I1(w11), .Z(s2));   //: @(650,619) /sn:0 /R:3 /w:[ 13 5 1 ]
  modul2 g48 (.H(w21), .G(w21), .S(w3), .Sk(s3));   //: @(563, 474) /sz:(60, 46) /sn:0 /p:[ Ti0>11 Ti1>9 Ti2>1 Bo0<0 ]
  //: joint g43 (w21) @(660, 407) /w:[ -1 1 2 12 ]
  //: joint g73 (w4) @(239, 473) /w:[ -1 5 6 8 ]
  //: joint g62 (w19) @(417, 291) /w:[ -1 1 2 4 ]
  modul1 g29 (.Pi(w11), .Gi(w10), .Pk(w15), .Gk(w14), .Pki(w20), .Gki(w13));   //: @(434, 296) /sz:(107, 63) /sn:0 /p:[ Ti0>3 Ti1>3 Ti2>5 Ti3>0 Bo0<1 Bo1<0 ]
  //: joint g25 (y3) @(504, 68) /w:[ -1 1 2 4 ]
  //: IN g17 (x1) @(663,30) /sn:0 /R:3 /w:[ 0 ]
  //: joint g88 (w33) @(22, 609) /w:[ 2 -1 4 1 ]
  //: joint g63 (w25) @(460, 647) /w:[ 4 -1 3 6 ]
  _GGXOR2 #(8) g52 (.I0(w26), .I1(w31), .Z(w36));   //: @(161,345) /sn:0 /R:3 /w:[ 5 3 1 ]
  modul1 g42 (.Pi(w24), .Gi(w21), .Pk(w20), .Gk(w13), .Pki(w25), .Gki(w12));   //: @(436, 522) /sz:(107, 63) /sn:0 /p:[ Ti0>5 Ti1>7 Ti2>0 Ti3>1 Bo0<5 Bo1<9 ]
  //: joint g83 (w12) @(161, 626) /w:[ 4 -1 3 14 ]
  //: joint g74 (w16) @(250, 449) /w:[ 4 -1 3 6 ]
  //: joint g56 (w31) @(140, 240) /w:[ 2 1 -1 4 ]
  //: IN g14 (y6) @(235,29) /sn:0 /R:3 /w:[ 0 ]
  generacja g5 (.y(y5), .x(x5), .h(w23), .g(w22));   //: @(271, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>5 Bo0<5 Bo1<0 ]
  //: joint g47 (w10) @(571, 266) /w:[ 1 -1 2 4 ]
  //: joint g44 (w24) @(552, 444) /w:[ 2 4 1 -1 ]
  //: joint g79 (w38) @(213, 460) /w:[ 6 -1 5 12 ]
  //: joint g80 (w16) @(157, 449) /w:[ 2 -1 1 8 ]
  //: joint g36 (w2) @(764, 274) /w:[ -1 2 1 4 ]
  //: joint g24 (y2) @(609, 45) /w:[ 2 1 -1 4 ]
  //: IN g21 (x5) @(294,29) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g84 (s7) @(160,805) /sn:0 /R:3 /w:[ 1 ]
  modul1 g85 (.Gk(w32), .Pk(w33), .Gi(w12), .Pi(w25), .Gki(c8), .Pki(w28));   //: @(-23, 693) /sz:(107, 63) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Bo0<0 Bo1<0 ]
  //: OUT g41 (s2) @(656,693) /sn:0 /R:3 /w:[ 0 ]
  //: IN g23 (x7) @(102,27) /sn:0 /R:3 /w:[ 0 ]
  //: joint g60 (w38) @(104, 460) /w:[ 2 1 -1 16 ]
  //: joint g54 (w23) @(330, 260) /w:[ 2 4 -1 1 ]
  //: joint g40 (w11) @(613, 280) /w:[ -1 1 2 4 ]
  //: joint g81 (w38) @(178, 460) /w:[ 4 -1 3 14 ]
  _GGAND2 #(6) g70 (.I0(w4), .I1(w38), .Z(w35));   //: @(218,508) /sn:0 /R:3 /w:[ 7 13 0 ]
  //: joint g46 (w15) @(508, 248) /w:[ 2 1 -1 4 ]
  _GGXOR2 #(8) g45 (.I0(w10), .I1(w15), .Z(w3));   //: @(567,361) /sn:0 /R:3 /w:[ 5 3 0 ]
  _GGXOR2 #(8) g35 (.I0(w2), .I1(w7), .Z(s1));   //: @(762,603) /sn:0 /R:3 /w:[ 5 3 0 ]
  //: joint g26 (x5) @(286, 49) /w:[ 1 2 -1 4 ]
  //: IN g22 (x6) @(203,31) /sn:0 /R:3 /w:[ 0 ]
  generacja g0 (.y(y0), .x(x0), .h(s0), .g(w2));   //: @(740, 78) /sz:(82, 91) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<3 ]
  //: joint g66 (w19) @(455, 665) /w:[ -1 5 6 8 ]
  modul2 g82 (.S(w39), .G(w12), .H(w35), .Sk(s7));   //: @(128, 697) /sz:(60, 46) /sn:0 /p:[ Ti0>0 Ti1>15 Ti2>1 Bo0<0 ]
  //: IN g18 (x2) @(564,30) /sn:0 /R:3 /w:[ 0 ]
  //: IN g12 (y4) @(412,28) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g33 (s0) @(809,620) /sn:0 /R:3 /w:[ 3 ]
  modul1 g30 (.Pi(s0), .Gi(w2), .Pk(w7), .Gk(w6), .Pki(w24), .Gki(w21));   //: @(630, 307) /sz:(107, 63) /sn:0 /p:[ Ti0>5 Ti1>0 Ti2>9 Ti3>5 Bo0<3 Bo1<0 ]
  //: joint g49 (w21) @(594, 407) /w:[ 5 -1 6 8 ]

endmodule
//: /netlistEnd

//: /netlistBegin modul2
module modul2(H, G, Sk, S);
//: interface  /sz:(60, 46) /bd:[ Ti0>S(12/60) Ti1>G(31/60) Ti2>H(51/60) Bo0<Sk(28/60) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
output Sk;    //: /sn:0 {0}(355,245)(355,306)(356,306)(356,313){1}
input G;    //: /sn:0 {0}(374,110)(374,152)(391,152){1}
//: {2}(393,150)(393,145){3}
//: {4}(393,154)(393,162){5}
input H;    //: /sn:0 {0}(395,138)(400,138){1}
//: {2}(404,138)(415,138)(415,110){3}
//: {4}(402,140)(402,150)(398,150)(398,162){5}
input S;    //: /sn:0 {0}(336,106)(336,209)(353,209)(353,224){1}
wire w2;    //: /sn:0 {0}(395,183)(395,209)(358,209)(358,224){1}
//: enddecls

  _GGXOR2 #(8) g4 (.I0(w2), .I1(S), .Z(Sk));   //: @(355,235) /sn:0 /R:3 /w:[ 1 1 0 ]
  _GGAND2 #(6) g3 (.I0(H), .I1(G), .Z(w2));   //: @(395,173) /sn:0 /R:3 /w:[ 5 5 0 ]
  //: IN g2 (H) @(415,108) /sn:0 /R:3 /w:[ 3 ]
  //: IN g1 (G) @(374,108) /sn:0 /R:3 /w:[ 0 ]
  //: joint g6 (H) @(402, 138) /w:[ 2 -1 1 4 ]
  //: OUT g7 (Sk) @(356,310) /sn:0 /R:3 /w:[ 1 ]
  //: joint g5 (G) @(393, 152) /w:[ -1 2 1 4 ]
  //: IN g0 (S) @(336,104) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin modul1
module modul1(Pi, Gi, Pk, Pki, Gki, Gk);
//: interface  /sz:(107, 63) /bd:[ Ti0>Gk(16/107) Ti1>Pk(33/107) Ti2>Gi(75/107) Ti3>Pi(92/107) Bo0<Gki(30/107) Bo1<Pki(59/107) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input Pk;    //: /sn:0 {0}(212,119)(212,87){1}
//: {2}(214,85)(277,85)(277,119){3}
//: {4}(212,83)(212,63){5}
output Gki;    //: /sn:0 {0}(195,287)(195,220){1}
output Pki;    //: /sn:0 {0}(279,140)(279,286){1}
input Gi;    //: /sn:0 {0}(217,119)(217,111)(256,111)(256,63){1}
input Gk;    //: /sn:0 {0}(172,63)(172,182)(193,182)(193,199){1}
input Pi;    //: /sn:0 {0}(317,63)(317,103)(282,103)(282,119){1}
wire w2;    //: /sn:0 {0}(214,140)(214,184)(198,184)(198,199){1}
//: enddecls

  //: joint g8 (Pk) @(212, 85) /w:[ 2 4 -1 1 ]
  _GGAND2 #(6) g4 (.I0(Gi), .I1(Pk), .Z(w2));   //: @(214,130) /sn:0 /R:3 /w:[ 0 0 0 ]
  //: IN g3 (Pi) @(317,61) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (Gi) @(256,61) /sn:0 /R:3 /w:[ 1 ]
  //: IN g1 (Pk) @(212,61) /sn:0 /R:3 /w:[ 5 ]
  _GGOR2 #(6) g6 (.I0(w2), .I1(Gk), .Z(Gki));   //: @(195,210) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: OUT g9 (Pki) @(279,283) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g7 (Gki) @(195,284) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g5 (.I0(Pi), .I1(Pk), .Z(Pki));   //: @(279,130) /sn:0 /R:3 /w:[ 1 3 0 ]
  //: IN g0 (Gk) @(172,61) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

